    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine �χ`    Q��!    q/0081;5ec14319;Chrome;AF5055D5-365C-4AF6-B333-CFCAC3BD1476 