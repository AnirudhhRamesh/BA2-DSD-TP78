    Mac OS X            	   2  >     p                                      ATTR      p   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     4   <  com.apple.quarantine ;ɇ`    �L:     ��6�JC�O-���C                                                      q/0081;5ea7e9e2;Chrome;9EEE266E-0C19-4EC9-ACF0-8993C160B99D 