    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine cƂ`    P�
(    q/0081;5eccebb3;Chrome;4B1A9969-1BC3-4416-8722-E0B0FD1F823E 